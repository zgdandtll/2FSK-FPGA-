library verilog;
use verilog.vl_types.all;
entity tb_tiaozhi is
end tb_tiaozhi;
