library verilog;
use verilog.vl_types.all;
entity jietiao_tb is
end jietiao_tb;
